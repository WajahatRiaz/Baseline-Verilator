`ifndef _HEADER_GUARD_
`define _HEADER_GUARD

`define MAX_DELAY #5
`define MIN_DELAY #2
`define CLOCK_HPERIOD #3
`define TIMEOUT #100
`endif